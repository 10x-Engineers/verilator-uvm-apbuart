`include "./../uvm_tb/apbinterface.sv" 
`include "./../uvm_tb/uartinterface.sv"
`include "./../uvm_tb/apb_transaction.sv" 
`include "./../uvm_tb/uart_transaction.sv" 
`include "./../uvm_tb/uart_config.sv"
`include "./../uvm_tb/apb_config.sv"
`include "./../uvm_tb/apb_sequencer.sv" 
`include "./../uvm_tb/uart_sequencer.sv"
`include "./../uvm_tb/apb_sequence.sv"
`include "./../uvm_tb/uart_sequence.sv" 
`include "./../uvm_tb/apbuart_vsequencer.sv" 
`include "./../uvm_tb/apbuart_vseq_base.sv" 
`include "./../uvm_tb/apb_driver.sv"
`include "./../uvm_tb/uart_driver.sv" 
`include "./../uvm_tb/apb_monitor.sv" 
`include "./../uvm_tb/uart_monitor.sv" 
`include "./../uvm_tb/apb_agent.sv"
`include "./../uvm_tb/uart_agent.sv" 
`include "./../uvm_tb/apbuart_scoreboard.sv" 
`include "./../uvm_tb/apbuart_environment.sv" 
`include "./../uvm_tb/apbuart_base_test.sv" 
`include "./../uvm_tb/apbuart_property.sv" 
`include "./../uvm_tb/apbuart_config_test.sv" 
`include "./../uvm_tb/apbuart_data_compare_test.sv" 
`include "./../uvm_tb/apbuart_parity_error_test.sv" 
`include "./../uvm_tb/apbuart_frame_error_test.sv" 
`include "./../uvm_tb/apbuart_free_error_test.sv" 
`include "./../uvm_tb/apbuart_rec_drv_test.sv"
`include "./../uvm_tb/apbuart_rec_readreg_test.sv"
